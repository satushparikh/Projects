library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;	 
use ieee.std_logic_unsigned.all;

-- since The Memory is asynchronous read, there is no read signal, but you can use it based on your preference.
-- this memory gives 16 Bit data in one clock cycle, so edit the file to your requirement.

entity Memory_Data is 
	port (address,Mem_datain: in std_logic_vector(15 downto 0); clk,Mem_wr: in std_logic;
				Mem_dataout: out std_logic_vector(15 downto 0));
end entity;

architecture ARC of Memory_Data is 
type regarray is array(65535 downto 0) of std_logic_vector(15 downto 0);   -- defining a new type
signal Memory: regarray:=(
   0 => x"0000" ,
   1 => x"0001" ,
   2 => x"0002" ,
   3 => x"0003" ,
   4 => x"0004" ,
   5 => x"0005" ,
   6 => x"0006" ,
   7 => x"0007" ,
   8 => x"0008" ,
   9 => x"0009" ,
   10 => x"000a" ,
   11 => x"000b" ,
   12 => x"000c" ,
   13 => x"000d" ,
   14 => x"000e" ,
   15 => x"000f" ,
   16 => x"0010" ,
   17 => x"0011" ,
   18 => x"0012" ,
   19 => x"0013" ,
   20 => x"0014" ,
   21 => x"0015" ,
   22 => x"0016" ,
   23 => x"0017" ,
   24 => x"0018" ,
   25 => x"0019" ,
   26 => x"001a" ,
   27 => x"001b" ,
   28 => x"001c" ,
   29 => x"001d" ,
   30 => x"001e" ,
   31 => x"001f" ,
   32 => x"0020" ,
   33 => x"0021" ,
   34 => x"0022" ,
   35 => x"0023" ,
   36 => x"0024" ,
   37 => x"0025" ,
   38 => x"0026" ,
   39 => x"0027" ,
   40 => x"0028" ,
   41 => x"0029" ,
   42 => x"002a" ,
   43 => x"002b" ,
   44 => x"002c" ,
   45 => x"002d" ,
   46 => x"002e" ,
   47 => x"002f" ,
   48 => x"0030" ,
   49 => x"0031" ,
   50 => x"0032" ,
   51 => x"0033" ,
   52 => x"0034" ,
   53 => x"0035" ,
   54 => x"0036" ,
   55 => x"0037" ,
   56 => x"0038" ,
   57 => x"0039" ,
   58 => x"003a" ,
   59 => x"003b" ,
   60 => x"003c" ,
   61 => x"003d" ,
   62 => x"003e" ,
   63 => x"003f" ,
   64 => x"0040" ,
   65 => x"0041" ,
   66 => x"0042" ,
   67 => x"0043" ,
   68 => x"0044" ,
   69 => x"0045" ,
   70 => x"0046" ,
   71 => x"0047" ,
   72 => x"0048" ,
   73 => x"0049" ,
   74 => x"004a" ,
   75 => x"004b" ,
   76 => x"004c" ,
   77 => x"004d" ,
   78 => x"004e" ,
   79 => x"004f" ,
   80 => x"0050" ,
   81 => x"0051" ,
   82 => x"0052" ,
   83 => x"0053" ,
   84 => x"0054" ,
   85 => x"0055" ,
   86 => x"0056" ,
   87 => x"0057" ,
   88 => x"0058" ,
   89 => x"0059" ,
   90 => x"005a" ,
   91 => x"005b" ,
   92 => x"005c" ,
   93 => x"005d" ,
   94 => x"005e" ,
   95 => x"005f" ,
   96 => x"0060" ,
   97 => x"0061" ,
   98 => x"0062" ,
   99 => x"0063" ,
   100 => x"0064" ,
   101 => x"0065" ,
   102 => x"0066" ,
   103 => x"0067" ,
   104 => x"0068" ,
   105 => x"0069" ,
   106 => x"006a" ,
   107 => x"006b" ,
   108 => x"006c" ,
   109 => x"006d" ,
   110 => x"006e" ,
   111 => x"006f" ,
   112 => x"0070" ,
   113 => x"0071" ,
   114 => x"0072" ,
   115 => x"0073" ,
   116 => x"0074" ,
   117 => x"0075" ,
   118 => x"0076" ,
   119 => x"0077" ,
   120 => x"0078" ,
   121 => x"0079" ,
   122 => x"007a" ,
   123 => x"007b" ,
   124 => x"007c" ,
   125 => x"007d" ,
   126 => x"007e" ,
   127 => x"007f" ,
   128 => x"0080" ,
   129 => x"0081" ,
   130 => x"0082" ,
   131 => x"0083" ,
   132 => x"0084" ,
   133 => x"0085" ,
   134 => x"0086" ,
   135 => x"0087" ,
   136 => x"0088" ,
   137 => x"0089" ,
   138 => x"008a" ,
   139 => x"008b" ,
   140 => x"008c" ,
   141 => x"008d" ,
   142 => x"008e" ,
   143 => x"008f" ,
   144 => x"0090" ,
   145 => x"0091" ,
   146 => x"0092" ,
   147 => x"0093" ,
   148 => x"0094" ,
   149 => x"0095" ,
   150 => x"0096" ,
   151 => x"0097" ,
   152 => x"0098" ,
   153 => x"0099" ,
   154 => x"009a" ,
   155 => x"009b" ,
   156 => x"009c" ,
   157 => x"009d" ,
   158 => x"009e" ,
   159 => x"009f" ,
   160 => x"00a0" ,
   161 => x"00a1" ,
   162 => x"00a2" ,
   163 => x"00a3" ,
   164 => x"00a4" ,
   165 => x"00a5" ,
   166 => x"00a6" ,
   167 => x"00a7" ,
   168 => x"00a8" ,
   169 => x"00a9" ,
   170 => x"00aa" ,
   171 => x"00ab" ,
   172 => x"00ac" ,
   173 => x"00ad" ,
   174 => x"00ae" ,
   175 => x"00af" ,
   176 => x"00b0" ,
   177 => x"00b1" ,
   178 => x"00b2" ,
   179 => x"00b3" ,
   180 => x"00b4" ,
   181 => x"00b5" ,
   182 => x"00b6" ,
   183 => x"00b7" ,
   184 => x"00b8" ,
   185 => x"00b9" ,
   186 => x"00ba" ,
   187 => x"00bb" ,
   188 => x"00bc" ,
   189 => x"00bd" ,
   190 => x"00be" ,
   191 => x"00bf" ,
   192 => x"00c0" ,
   193 => x"00c1" ,
   194 => x"00c2" ,
   195 => x"00c3" ,
   196 => x"00c4" ,
   197 => x"00c5" ,
   198 => x"00c6" ,
   199 => x"00c7" ,
   200 => x"00c8" ,
   201 => x"00c9" ,
   202 => x"00ca" ,
   203 => x"00cb" ,
   204 => x"00cc" ,
   205 => x"00cd" ,
   206 => x"00ce" ,
   207 => x"00cf" ,
   208 => x"00d0" ,
   209 => x"00d1" ,
   210 => x"00d2" ,
   211 => x"00d3" ,
   212 => x"00d4" ,
   213 => x"00d5" ,
   214 => x"00d6" ,
   215 => x"00d7" ,
   216 => x"00d8" ,
   217 => x"00d9" ,
   218 => x"00da" ,
   219 => x"00db" ,
   220 => x"00dc" ,
   221 => x"00dd" ,
   222 => x"00de" ,
   223 => x"00df" ,
   224 => x"00e0" ,
   225 => x"00e1" ,
   226 => x"00e2" ,
   227 => x"00e3" ,
   228 => x"00e4" ,
   229 => x"00e5" ,
   230 => x"00e6" ,
   231 => x"00e7" ,
   232 => x"00e8" ,
   233 => x"00e9" ,
   234 => x"00ea" ,
   235 => x"00eb" ,
   236 => x"00ec" ,
   237 => x"00ed" ,
   238 => x"00ee" ,
   239 => x"00ef" ,
   240 => x"00f0" ,
   241 => x"00f1" ,
   242 => x"00f2" ,
   243 => x"00f3" ,
   244 => x"00f4" ,
   245 => x"00f5" ,
   246 => x"00f6" ,
   247 => x"00f7" ,
   248 => x"00f8" ,
   249 => x"00f9" ,
   250 => x"00fa" ,
   251 => x"00fb" ,
   252 => x"00fc" ,
   253 => x"00fd" ,
   254 => x"00fe" ,
   255 => x"00ff" ,
   256 => x"0100" ,
   257 => x"0101" ,
   258 => x"0102" ,
   259 => x"0103" ,
   260 => x"0104" ,
   261 => x"0105" ,
   262 => x"0106" ,
   263 => x"0107" ,
   264 => x"0108" ,
   265 => x"0109" ,
   266 => x"010a" ,
   267 => x"010b" ,
   268 => x"010c" ,
   269 => x"010d" ,
   270 => x"010e" ,
   271 => x"010f" ,
   272 => x"0110" ,
   273 => x"0111" ,
   274 => x"0112" ,
   275 => x"0113" ,
   276 => x"0114" ,
   277 => x"0115" ,
   278 => x"0116" ,
   279 => x"0117" ,
   280 => x"0118" ,
   281 => x"0119" ,
   282 => x"011a" ,
   283 => x"011b" ,
   284 => x"011c" ,
   285 => x"011d" ,
   286 => x"011e" ,
   287 => x"011f" ,
   288 => x"0120" ,
   289 => x"0121" ,
   290 => x"0122" ,
   291 => x"0123" ,
   292 => x"0124" ,
   293 => x"0125" ,
   294 => x"0126" ,
   295 => x"0127" ,
   296 => x"0128" ,
   297 => x"0129" ,
   298 => x"012a" ,
   299 => x"012b" ,
   300 => x"012c" ,
   301 => x"012d" ,
   302 => x"012e" ,
   303 => x"012f" ,
   304 => x"0130" ,
   305 => x"0131" ,
   306 => x"0132" ,
   307 => x"0133" ,
   308 => x"0134" ,
   309 => x"0135" ,
   310 => x"0136" ,
   311 => x"0137" ,
   312 => x"0138" ,
   313 => x"0139" ,
   314 => x"013a" ,
   315 => x"013b" ,
   316 => x"013c" ,
   317 => x"013d" ,
   318 => x"013e" ,
   319 => x"013f" ,
   320 => x"0140" ,
   321 => x"0141" ,
   322 => x"0142" ,
   323 => x"0143" ,
   324 => x"0144" ,
   325 => x"0145" ,
   326 => x"0146" ,
   327 => x"0147" ,
   328 => x"0148" ,
   329 => x"0149" ,
   330 => x"014a" ,
   331 => x"014b" ,
   332 => x"014c" ,
   333 => x"014d" ,
   334 => x"014e" ,
   335 => x"014f" ,
   336 => x"0150" ,
   337 => x"0151" ,
   338 => x"0152" ,
   339 => x"0153" ,
   340 => x"0154" ,
   341 => x"0155" ,
   342 => x"0156" ,
   343 => x"0157" ,
   344 => x"0158" ,
   345 => x"0159" ,
   346 => x"015a" ,
   347 => x"015b" ,
   348 => x"015c" ,
   349 => x"015d" ,
   350 => x"015e" ,
   351 => x"015f" ,
   352 => x"0160" ,
   353 => x"0161" ,
   354 => x"0162" ,
   355 => x"0163" ,
   356 => x"0164" ,
   357 => x"0165" ,
   358 => x"0166" ,
   359 => x"0167" ,
   360 => x"0168" ,
   361 => x"0169" ,
   362 => x"016a" ,
   363 => x"016b" ,
   364 => x"016c" ,
   365 => x"016d" ,
   366 => x"016e" ,
   367 => x"016f" ,
   368 => x"0170" ,
   369 => x"0171" ,
   370 => x"0172" ,
   371 => x"0173" ,
   372 => x"0174" ,
   373 => x"0175" ,
   374 => x"0176" ,
   375 => x"0177" ,
   376 => x"0178" ,
   377 => x"0179" ,
   378 => x"017a" ,
   379 => x"017b" ,
   380 => x"017c" ,
   381 => x"017d" ,
   382 => x"017e" ,
   383 => x"017f" ,
   384 => x"0180" ,
   385 => x"0181" ,
   386 => x"0182" ,
   387 => x"0183" ,
   388 => x"0184" ,
   389 => x"0185" ,
   390 => x"0186" ,
   391 => x"0187" ,
   392 => x"0188" ,
   393 => x"0189" ,
   394 => x"018a" ,
   395 => x"018b" ,
   396 => x"018c" ,
   397 => x"018d" ,
   398 => x"018e" ,
   399 => x"018f" ,
   400 => x"0190" ,
   401 => x"0191" ,
   402 => x"0192" ,
   403 => x"0193" ,
   404 => x"0194" ,
   405 => x"0195" ,
   406 => x"0196" ,
   407 => x"0197" ,
   408 => x"0198" ,
   409 => x"0199" ,
   410 => x"019a" ,
   411 => x"019b" ,
   412 => x"019c" ,
   413 => x"019d" ,
   414 => x"019e" ,
   415 => x"019f" ,
   416 => x"01a0" ,
   417 => x"01a1" ,
   418 => x"01a2" ,
   419 => x"01a3" ,
   420 => x"01a4" ,
   421 => x"01a5" ,
   422 => x"01a6" ,
   423 => x"01a7" ,
   424 => x"01a8" ,
   425 => x"01a9" ,
   426 => x"01aa" ,
   427 => x"01ab" ,
   428 => x"01ac" ,
   429 => x"01ad" ,
   430 => x"01ae" ,
   431 => x"01af" ,
   432 => x"01b0" ,
   433 => x"01b1" ,
   434 => x"01b2" ,
   435 => x"01b3" ,
   436 => x"01b4" ,
   437 => x"01b5" ,
   438 => x"01b6" ,
   439 => x"01b7" ,
   440 => x"01b8" ,
   441 => x"01b9" ,
   442 => x"01ba" ,
   443 => x"01bb" ,
   444 => x"01bc" ,
   445 => x"01bd" ,
   446 => x"01be" ,
   447 => x"01bf" ,
   448 => x"01c0" ,
   449 => x"01c1" ,
   450 => x"01c2" ,
   451 => x"01c3" ,
   452 => x"01c4" ,
   453 => x"01c5" ,
   454 => x"01c6" ,
   455 => x"01c7" ,
   456 => x"01c8" ,
   457 => x"01c9" ,
   458 => x"01ca" ,
   459 => x"01cb" ,
   460 => x"01cc" ,
   461 => x"01cd" ,
   462 => x"01ce" ,
   463 => x"01cf" ,
   464 => x"01d0" ,
   465 => x"01d1" ,
   466 => x"01d2" ,
   467 => x"01d3" ,
   468 => x"01d4" ,
   469 => x"01d5" ,
   470 => x"01d6" ,
   471 => x"01d7" ,
   472 => x"01d8" ,
   473 => x"01d9" ,
   474 => x"01da" ,
   475 => x"01db" ,
   476 => x"01dc" ,
   477 => x"01dd" ,
   478 => x"01de" ,
   479 => x"01df" ,
   480 => x"01e0" ,
   481 => x"01e1" ,
   482 => x"01e2" ,
   483 => x"01e3" ,
   484 => x"01e4" ,
   485 => x"01e5" ,
   486 => x"01e6" ,
   487 => x"01e7" ,
   488 => x"01e8" ,
   489 => x"01e9" ,
   490 => x"01ea" ,
   491 => x"01eb" ,
   492 => x"01ec" ,
   493 => x"01ed" ,
   494 => x"01ee" ,
   495 => x"01ef" ,
   496 => x"01f0" ,
   497 => x"01f1" ,
   498 => x"01f2" ,
   499 => x"01f3" ,
   500 => x"01f4" ,
   501 => x"01f5" ,
   502 => x"01f6" ,
   503 => x"01f7" ,
   504 => x"01f8" ,
   505 => x"01f9" ,
   506 => x"01fa" ,
   507 => x"01fb" ,
   508 => x"01fc" ,
   509 => x"01fd" ,
   510 => x"01fe" ,
   511 => x"01ff" ,
   512 => x"0200" ,
   513 => x"0201" ,
   514 => x"0202" ,
   515 => x"0203" ,
   516 => x"0204" ,
   517 => x"0205" ,
   518 => x"0206" ,
   519 => x"0207" ,
   520 => x"0208" ,
   521 => x"0209" ,
   522 => x"020a" ,
   523 => x"020b" ,
   524 => x"020c" ,
   525 => x"020d" ,
   526 => x"020e" ,
   527 => x"020f" ,
   528 => x"0210" ,
   529 => x"0211" ,
   530 => x"0212" ,
   531 => x"0213" ,
   532 => x"0214" ,
   533 => x"0215" ,
   534 => x"0216" ,
   535 => x"0217" ,
   536 => x"0218" ,
   537 => x"0219" ,
   538 => x"021a" ,
   539 => x"021b" ,
   540 => x"021c" ,
   541 => x"021d" ,
   542 => x"021e" ,
   543 => x"021f" ,
   544 => x"0220" ,
   545 => x"0221" ,
   546 => x"0222" ,
   547 => x"0223" ,
   548 => x"0224" ,
   549 => x"0225" ,
   550 => x"0226" ,
   551 => x"0227" ,
   552 => x"0228" ,
   553 => x"0229" ,
   554 => x"022a" ,
   555 => x"022b" ,
   556 => x"022c" ,
   557 => x"022d" ,
   558 => x"022e" ,
   559 => x"022f" ,
   560 => x"0230" ,
   561 => x"0231" ,
   562 => x"0232" ,
   563 => x"0233" ,
   564 => x"0234" ,
   565 => x"0235" ,
   566 => x"0236" ,
   567 => x"0237" ,
   568 => x"0238" ,
   569 => x"0239" ,
   570 => x"023a" ,
   571 => x"023b" ,
   572 => x"023c" ,
   573 => x"023d" ,
   574 => x"023e" ,
   575 => x"023f" ,
   576 => x"0240" ,
   577 => x"0241" ,
   578 => x"0242" ,
   579 => x"0243" ,
   580 => x"0244" ,
   581 => x"0245" ,
   582 => x"0246" ,
   583 => x"0247" ,
   584 => x"0248" ,
   585 => x"0249" ,
   586 => x"024a" ,
   587 => x"024b" ,
   588 => x"024c" ,
   589 => x"024d" ,
   590 => x"024e" ,
   591 => x"024f" ,
   592 => x"0250" ,
   593 => x"0251" ,
   594 => x"0252" ,
   595 => x"0253" ,
   596 => x"0254" ,
   597 => x"0255" ,
   598 => x"0256" ,
   599 => x"0257" ,
   600 => x"0258" ,
   601 => x"0259" ,
   602 => x"025a" ,
   603 => x"025b" ,
   604 => x"025c" ,
   605 => x"025d" ,
   606 => x"025e" ,
   607 => x"025f" ,
   608 => x"0260" ,
   609 => x"0261" ,
   610 => x"0262" ,
   611 => x"0263" ,
   612 => x"0264" ,
   613 => x"0265" ,
   614 => x"0266" ,
   615 => x"0267" ,
   616 => x"0268" ,
   617 => x"0269" ,
   618 => x"026a" ,
   619 => x"026b" ,
   620 => x"026c" ,
   621 => x"026d" ,
   622 => x"026e" ,
   623 => x"026f" ,
   624 => x"0270" ,
   625 => x"0271" ,
   626 => x"0272" ,
   627 => x"0273" ,
   628 => x"0274" ,
   629 => x"0275" ,
   630 => x"0276" ,
   631 => x"0277" ,
   632 => x"0278" ,
   633 => x"0279" ,
   634 => x"027a" ,
   635 => x"027b" ,
   636 => x"027c" ,
   637 => x"027d" ,
   638 => x"027e" ,
   639 => x"027f" ,
   640 => x"0280" ,
   641 => x"0281" ,
   642 => x"0282" ,
   643 => x"0283" ,
   644 => x"0284" ,
   645 => x"0285" ,
   646 => x"0286" ,
   647 => x"0287" ,
   648 => x"0288" ,
   649 => x"0289" ,
   650 => x"028a" ,
   651 => x"028b" ,
   652 => x"028c" ,
   653 => x"028d" ,
   654 => x"028e" ,
   655 => x"028f" ,
   656 => x"0290" ,
   657 => x"0291" ,
   658 => x"0292" ,
   659 => x"0293" ,
   660 => x"0294" ,
   661 => x"0295" ,
   662 => x"0296" ,
   663 => x"0297" ,
   664 => x"0298" ,
   665 => x"0299" ,
   666 => x"029a" ,
   667 => x"029b" ,
   668 => x"029c" ,
   669 => x"029d" ,
   670 => x"029e" ,
   671 => x"029f" ,
   672 => x"02a0" ,
   673 => x"02a1" ,
   674 => x"02a2" ,
   675 => x"02a3" ,
   676 => x"02a4" ,
   677 => x"02a5" ,
   678 => x"02a6" ,
   679 => x"02a7" ,
   680 => x"02a8" ,
   681 => x"02a9" ,
   682 => x"02aa" ,
   683 => x"02ab" ,
   684 => x"02ac" ,
   685 => x"02ad" ,
   686 => x"02ae" ,
   687 => x"02af" ,
   688 => x"02b0" ,
   689 => x"02b1" ,
   690 => x"02b2" ,
   691 => x"02b3" ,
   692 => x"02b4" ,
   693 => x"02b5" ,
   694 => x"02b6" ,
   695 => x"02b7" ,
   696 => x"02b8" ,
   697 => x"02b9" ,
   698 => x"02ba" ,
   699 => x"02bb" ,
   700 => x"02bc" ,
   701 => x"02bd" ,
   702 => x"02be" ,
   703 => x"02bf" ,
   704 => x"02c0" ,
   705 => x"02c1" ,
   706 => x"02c2" ,
   707 => x"02c3" ,
   708 => x"02c4" ,
   709 => x"02c5" ,
   710 => x"02c6" ,
   711 => x"02c7" ,
   712 => x"02c8" ,
   713 => x"02c9" ,
   714 => x"02ca" ,
   715 => x"02cb" ,
   716 => x"02cc" ,
   717 => x"02cd" ,
   718 => x"02ce" ,
   719 => x"02cf" ,
   720 => x"02d0" ,
   721 => x"02d1" ,
   722 => x"02d2" ,
   723 => x"02d3" ,
   724 => x"02d4" ,
   725 => x"02d5" ,
   726 => x"02d6" ,
   727 => x"02d7" ,
   728 => x"02d8" ,
   729 => x"02d9" ,
   730 => x"02da" ,
   731 => x"02db" ,
   732 => x"02dc" ,
   733 => x"02dd" ,
   734 => x"02de" ,
   735 => x"02df" ,
   736 => x"02e0" ,
   737 => x"02e1" ,
   738 => x"02e2" ,
   739 => x"02e3" ,
   740 => x"02e4" ,
   741 => x"02e5" ,
   742 => x"02e6" ,
   743 => x"02e7" ,
   744 => x"02e8" ,
   745 => x"02e9" ,
   746 => x"02ea" ,
   747 => x"02eb" ,
   748 => x"02ec" ,
   749 => x"02ed" ,
   750 => x"02ee" ,
   751 => x"02ef" ,
   752 => x"02f0" ,
   753 => x"02f1" ,
   754 => x"02f2" ,
   755 => x"02f3" ,
   756 => x"02f4" ,
   757 => x"02f5" ,
   758 => x"02f6" ,
   759 => x"02f7" ,
   760 => x"02f8" ,
   761 => x"02f9" ,
   762 => x"02fa" ,
   763 => x"02fb" ,
   764 => x"02fc" ,
   765 => x"02fd" ,
   766 => x"02fe" ,
   767 => x"02ff" ,
   768 => x"0300" ,
   769 => x"0301" ,
   770 => x"0302" ,
   771 => x"0303" ,
   772 => x"0304" ,
   773 => x"0305" ,
   774 => x"0306" ,
   775 => x"0307" ,
   776 => x"0308" ,
   777 => x"0309" ,
   778 => x"030a" ,
   779 => x"030b" ,
   780 => x"030c" ,
   781 => x"030d" ,
   782 => x"030e" ,
   783 => x"030f" ,
   784 => x"0310" ,
   785 => x"0311" ,
   786 => x"0312" ,
   787 => x"0313" ,
   788 => x"0314" ,
   789 => x"0315" ,
   790 => x"0316" ,
   791 => x"0317" ,
   792 => x"0318" ,
   793 => x"0319" ,
   794 => x"031a" ,
   795 => x"031b" ,
   796 => x"031c" ,
   797 => x"031d" ,
   798 => x"031e" ,
   799 => x"031f" ,
   800 => x"0320" ,
   801 => x"0321" ,
   802 => x"0322" ,
   803 => x"0323" ,
   804 => x"0324" ,
   805 => x"0325" ,
   806 => x"0326" ,
   807 => x"0327" ,
   808 => x"0328" ,
   809 => x"0329" ,
   810 => x"032a" ,
   811 => x"032b" ,
   812 => x"032c" ,
   813 => x"032d" ,
   814 => x"032e" ,
   815 => x"032f" ,
   816 => x"0330" ,
   817 => x"0331" ,
   818 => x"0332" ,
   819 => x"0333" ,
   820 => x"0334" ,
   821 => x"0335" ,
   822 => x"0336" ,
   823 => x"0337" ,
   824 => x"0338" ,
   825 => x"0339" ,
   826 => x"033a" ,
   827 => x"033b" ,
   828 => x"033c" ,
   829 => x"033d" ,
   830 => x"033e" ,
   831 => x"033f" ,
   832 => x"0340" ,
   833 => x"0341" ,
   834 => x"0342" ,
   835 => x"0343" ,
   836 => x"0344" ,
   837 => x"0345" ,
   838 => x"0346" ,
   839 => x"0347" ,
   840 => x"0348" ,
   841 => x"0349" ,
   842 => x"034a" ,
   843 => x"034b" ,
   844 => x"034c" ,
   845 => x"034d" ,
   846 => x"034e" ,
   847 => x"034f" ,
   848 => x"0350" ,
   849 => x"0351" ,
   850 => x"0352" ,
   851 => x"0353" ,
   852 => x"0354" ,
   853 => x"0355" ,
   854 => x"0356" ,
   855 => x"0357" ,
   856 => x"0358" ,
   857 => x"0359" ,
   858 => x"035a" ,
   859 => x"035b" ,
   860 => x"035c" ,
   861 => x"035d" ,
   862 => x"035e" ,
   863 => x"035f" ,
   864 => x"0360" ,
   865 => x"0361" ,
   866 => x"0362" ,
   867 => x"0363" ,
   868 => x"0364" ,
   869 => x"0365" ,
   870 => x"0366" ,
   871 => x"0367" ,
   872 => x"0368" ,
   873 => x"0369" ,
   874 => x"036a" ,
   875 => x"036b" ,
   876 => x"036c" ,
   877 => x"036d" ,
   878 => x"036e" ,
   879 => x"036f" ,
   880 => x"0370" ,
   881 => x"0371" ,
   882 => x"0372" ,
   883 => x"0373" ,
   884 => x"0374" ,
   885 => x"0375" ,
   886 => x"0376" ,
   887 => x"0377" ,
   888 => x"0378" ,
   889 => x"0379" ,
   890 => x"037a" ,
   891 => x"037b" ,
   892 => x"037c" ,
   893 => x"037d" ,
   894 => x"037e" ,
   895 => x"037f" ,
   896 => x"0380" ,
   897 => x"0381" ,
   898 => x"0382" ,
   899 => x"0383" ,
   900 => x"0384" ,
   901 => x"0385" ,
   902 => x"0386" ,
   903 => x"0387" ,
   904 => x"0388" ,
   905 => x"0389" ,
   906 => x"038a" ,
   907 => x"038b" ,
   908 => x"038c" ,
   909 => x"038d" ,
   910 => x"038e" ,
   911 => x"038f" ,
   912 => x"0390" ,
   913 => x"0391" ,
   914 => x"0392" ,
   915 => x"0393" ,
   916 => x"0394" ,
   917 => x"0395" ,
   918 => x"0396" ,
   919 => x"0397" ,
   920 => x"0398" ,
   921 => x"0399" ,
   922 => x"039a" ,
   923 => x"039b" ,
   924 => x"039c" ,
   925 => x"039d" ,
   926 => x"039e" ,
   927 => x"039f" ,
   928 => x"03a0" ,
   929 => x"03a1" ,
   930 => x"03a2" ,
   931 => x"03a3" ,
   932 => x"03a4" ,
   933 => x"03a5" ,
   934 => x"03a6" ,
   935 => x"03a7" ,
   936 => x"03a8" ,
   937 => x"03a9" ,
   938 => x"03aa" ,
   939 => x"03ab" ,
   940 => x"03ac" ,
   941 => x"03ad" ,
   942 => x"03ae" ,
   943 => x"03af" ,
   944 => x"03b0" ,
   945 => x"03b1" ,
   946 => x"03b2" ,
   947 => x"03b3" ,
   948 => x"03b4" ,
   949 => x"03b5" ,
   950 => x"03b6" ,
   951 => x"03b7" ,
   952 => x"03b8" ,
   953 => x"03b9" ,
   954 => x"03ba" ,
   955 => x"03bb" ,
   956 => x"03bc" ,
   957 => x"03bd" ,
   958 => x"03be" ,
   959 => x"03bf" ,
   960 => x"03c0" ,
   961 => x"03c1" ,
   962 => x"03c2" ,
   963 => x"03c3" ,
   964 => x"03c4" ,
   965 => x"03c5" ,
   966 => x"03c6" ,
   967 => x"03c7" ,
   968 => x"03c8" ,
   969 => x"03c9" ,
   970 => x"03ca" ,
   971 => x"03cb" ,
   972 => x"03cc" ,
   973 => x"03cd" ,
   974 => x"03ce" ,
   975 => x"03cf" ,
   976 => x"03d0" ,
   977 => x"03d1" ,
   978 => x"03d2" ,
   979 => x"03d3" ,
   980 => x"03d4" ,
   981 => x"03d5" ,
   982 => x"03d6" ,
   983 => x"03d7" ,
   984 => x"03d8" ,
   985 => x"03d9" ,
   986 => x"03da" ,
   987 => x"03db" ,
   988 => x"03dc" ,
   989 => x"03dd" ,
   990 => x"03de" ,
   991 => x"03df" ,
   992 => x"03e0" ,
   993 => x"03e1" ,
   994 => x"03e2" ,
   995 => x"03e3" ,
   996 => x"03e4" ,
   997 => x"03e5" ,
   998 => x"03e6" ,
   999 => x"03e7" ,
   1000 => x"03e8" ,
   1001 => x"03e9" ,
   1002 => x"03ea" ,
   1003 => x"03eb" ,
   1004 => x"03ec" ,
   1005 => x"03ed" ,
   1006 => x"03ee" ,
   1007 => x"03ef" ,
   1008 => x"03f0" ,
   1009 => x"03f1" ,
   1010 => x"03f2" ,
   1011 => x"03f3" ,
   1012 => x"03f4" ,
   1013 => x"03f5" ,
   1014 => x"03f6" ,
   1015 => x"03f7" ,
   1016 => x"03f8" ,
   1017 => x"03f9" ,
   1018 => x"03fa" ,
   1019 => x"03fb" ,
   1020 => x"03fc" ,
   1021 => x"03fd" ,
   1022 => x"03fe" ,
   1023 => x"03ff" ,
    others => x"0000");

    begin
Mem_dataout <= Memory(conv_integer(address));
Mem_write:
process (Mem_wr,Mem_datain,address,clk)
	begin
	if(Mem_wr = '1') then
		if(rising_edge(clk)) then
			Memory(conv_integer(address)) <= Mem_datain;
		end if;
	end if;
	end process;
end ARC;
